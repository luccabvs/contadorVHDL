library IEEE;
use IEEE.std_logic_1164.all;
use ieee.numeric_std.all;

entity memoriaROM is
   generic (
          dataWidth: natural := 4;
          addrWidth: natural := 9
    );
   port (
          Endereco : in std_logic_vector (addrWidth-1 DOWNTO 0);
          Dado : out std_logic_vector (dataWidth-1 DOWNTO 0)
    );
end entity;

architecture assincrona of memoriaROM is

  type blocoMemoria is array(0 TO 2**addrWidth - 1) of std_logic_vector(dataWidth-1 DOWNTO 0);

  function initMemory
        return blocoMemoria is variable tmp : blocoMemoria := (others => (others => '0'));
		  
		  
  constant NOP  : std_logic_vector(3 downto 0) := "0000";
  constant LDA  : std_logic_vector(3 downto 0) := "0001";
  constant SOMA : std_logic_vector(3 downto 0) := "0010";
  constant SUB  : std_logic_vector(3 downto 0) := "0011";
  constant LDI  : std_logic_vector(3 downto 0) := "0100";
  constant STA  : std_logic_vector(3 downto 0) := "0101";
  constant JMP  : std_logic_vector(3 downto 0) := "0110";
  constant JEQ  : std_logic_vector(3 downto 0) := "0111";
  constant CEQ  : std_logic_vector(3 downto 0) := "1000";
  constant JSR  : std_logic_vector(3 downto 0) := "1001";
  constant RET  : std_logic_vector(3 downto 0) := "1010";

		  
		  
  begin
      -- Palavra de Controle = SelMUX, Habilita_A, Reset_A, Operacao_ULA
      -- Inicializa os endereços:

tmp(0) := NOP & '0' & x"00";	-- !Reset
tmp(1) := STA & '1' & x"FE";	-- STA @510                    	--Limpa leitura KEY1
tmp(2) := STA & '1' & x"FF";	-- STA @511                    	--Limpa leitura KEY0
tmp(3) := STA & '1' & x"FD";	-- STA @509                    	--Limpa leitura Reset    
tmp(4) := LDI & '0' & x"01";	-- LDI $1                      	--Carrega 1 no acumulador
tmp(5) := STA & '0' & x"3F";	-- STA @63                     	--Salva 1 no endereço 63 da RAM
tmp(6) := LDI & '0' & x"09";	-- LDI $9                      	--Carrega 9 no acumulador
tmp(7) := STA & '0' & x"13";	-- STA @19                     	--Salva 9 no endereço 19 da RAM
tmp(8) := LDI & '0' & x"0A";	-- LDI $10                     	--Carrega 10 no acumulador
tmp(9) := STA & '0' & x"14";	-- STA @20                     	--Salva 10 no endereço 20 da RAM
tmp(10) := LDI & '0' & x"0B";	-- LDI $11                     	--Carrega 11 no acumulador
tmp(11) := STA & '0' & x"15";	-- STA @21                     	--Salva 11 no endereço 21 da RAM
tmp(12) := LDI & '0' & x"0C";	-- LDI $12                     	--Carrega 12 no acumulador
tmp(13) := STA & '0' & x"16";	-- STA @22                     	--Salva 12 no endereço 22 da RAM
tmp(14) := LDI & '0' & x"0D";	-- LDI $13                     	--Carrega 13 no acumulador
tmp(15) := STA & '0' & x"17";	-- STA @23                     	--Salva 13 no endereço 23 da RAM
tmp(16) := LDI & '0' & x"0E";	-- LDI $14                     	--Carrega 14 no acumulador
tmp(17) := STA & '0' & x"18";	-- STA @24                     	--Salva 14 no endereço 24 da RAM
tmp(18) := LDI & '0' & x"0F";	-- LDI $15                     	--Carrega 15 no acumulador
tmp(19) := STA & '0' & x"19";	-- STA @25                     	--Salva 15 no endereço 25 da RAM
tmp(20) := LDI & '0' & x"00";	-- LDI $0                      	--Carrega 0 no acumulador
tmp(21) := STA & '0' & x"3E";	-- STA @62                     	--Salva 0 no endereço 62 da RAM
tmp(22) := STA & '1' & x"02";	-- STA @258                    	--Apaga o LED 9
tmp(23) := STA & '1' & x"01";	-- STA @257                    	--Apaga o LED 8
tmp(24) := STA & '1' & x"00";	-- STA @256                    	--Apaga o LED 7 a 0 
tmp(25) := STA & '1' & x"20";	-- STA @288                    	--Zera o HEX 0
tmp(26) := STA & '1' & x"21";	-- STA @289                    	--Zera o HEX 1
tmp(27) := STA & '1' & x"22";	-- STA @290                    	--Zera o HEX 2
tmp(28) := STA & '1' & x"23";	-- STA @291                    	--Zera o HEX 3
tmp(29) := STA & '1' & x"24";	-- STA @292                    	--Zera o HEX 4
tmp(30) := STA & '1' & x"25";	-- STA @293                    	--Zera o HEX 5
tmp(31) := STA & '0' & x"00";	-- STA @0                      	--Zera o endereço 0 da RAM (Limite das unidades)
tmp(32) := STA & '0' & x"01";	-- STA @1                      	--Zera o endereço 1 da RAM (Limite das dezenas)
tmp(33) := STA & '0' & x"02";	-- STA @2                      	--Zera o endereço 2 da RAM (Limite das centenas) 
tmp(34) := STA & '0' & x"03";	-- STA @3                      	--Zera o endereço 3 da RAM (Limite dos milhares) 
tmp(35) := STA & '0' & x"04";	-- STA @4                      	--Zera o endereço 4 da RAM (Limite das dezenas de milhares)
tmp(36) := STA & '0' & x"05";	-- STA @5                      	--Zera o endereço 5 da RAM (Limite das centenas de milhares) 
tmp(37) := STA & '0' & x"0A";	-- STA @10                     	--Zera o endereço 10 da RAM (Valor atual das unidades) 
tmp(38) := STA & '0' & x"0B";	-- STA @11                     	--Zera o endereço 11 da RAM (Valor atual das dezenas)
tmp(39) := STA & '0' & x"0C";	-- STA @12                     	--Zera o endereço 12 da RAM (Valor atual das centenas)
tmp(40) := STA & '0' & x"0D";	-- STA @13                     	--Zera o endereço 13 da RAM (Valor atual dos milhares)
tmp(41) := STA & '0' & x"0E";	-- STA @14                     	--Zera o endereço 14 da RAM (Valor atual das dezenas de milhares)
tmp(42) := STA & '0' & x"0F";	-- STA @15                     	--Zera o endereço 15 da RAM (Valor atual das centenas de milhares)
tmp(43) := NOP & '0' & x"00";	-- !Start
tmp(44) := LDA & '1' & x"61";	-- LDA @353                    	--Carrega o valor do KEY1 no acumulador
tmp(45) := CEQ & '0' & x"3F";	-- CEQ @63                     	--Compara o valor do KEY1 com 63 (1)
tmp(46) := JEQ & '0' & x"36";	-- JEQ @SetLim                 	--Se o valor do KEY1 for 1, vai para o label SetLim (Setar Limite)
tmp(47) := LDA & '1' & x"60";	-- LDA @352                    	--Carrega o valor do KEY0 no acumulador
tmp(48) := CEQ & '0' & x"3F";	-- CEQ @63                     	--Compara o valor do KEY0 com 63 (1)
tmp(49) := JEQ & '0' & x"ED";	-- JEQ @Incremento             	--Se o valor do KEY0 for 1, vai para o label Incremento (Incrementar)
tmp(50) := LDA & '1' & x"64";	-- LDA @356                    	--Carrega o valor do Reset no acumulador
tmp(51) := CEQ & '0' & x"3F";	-- CEQ @63                     	--Compara o valor do Reset com 63 (1)
tmp(52) := JEQ & '0' & x"00";	-- JEQ @Reset                  	--Se o valor do Reset for 1, vai para o label Reset (Reseta o programa)
tmp(53) := JMP & '0' & x"2B";	-- JMP @Start                  	--Se nenhum dos botoes forem clicados, vai para o label Start (Laco principal)
tmp(54) := NOP & '0' & x"00";	-- !SetLim
tmp(55) := STA & '1' & x"FE";	-- STA @510                    	--Limpa leitura KEY1
tmp(56) := LDA & '0' & x"00";	-- LDA @0                      	--Carrega o valor do endereço 0 da RAM no acumulador (Limite das unidades)
tmp(57) := STA & '1' & x"20";	-- STA @288                    	--Mostra o valor do acumulador HEX 0 (unidades)
tmp(58) := LDA & '0' & x"01";	-- LDA @1                      	--Carrega o valor do endereço 1 da RAM no acumulador (Limite das dezenas)
tmp(59) := STA & '1' & x"21";	-- STA @289                    	--Mostra o valor do acumulador HEX 1 (dezenas)
tmp(60) := LDA & '0' & x"02";	-- LDA @2                      	--Carrega o valor do endereço 2 da RAM no acumulador (Limite das centenas)
tmp(61) := STA & '1' & x"22";	-- STA @290                    	--Mostra o valor do acumulador HEX 2 (centenas)
tmp(62) := LDA & '0' & x"03";	-- LDA @3                      	--Carrega o valor do endereço 3 da RAM no acumulador (Limite dos milhares)
tmp(63) := STA & '1' & x"23";	-- STA @291                    	--Mostra o valor do acumulador HEX 3 (milhares)
tmp(64) := LDA & '0' & x"04";	-- LDA @4                      	--Carrega o valor do endereço 4 da RAM no acumulador (Limite das dezenas de milhares)
tmp(65) := STA & '1' & x"24";	-- STA @292                    	--Mostra o valor do acumulador HEX 4 (dezenas de milhares)
tmp(66) := LDA & '0' & x"05";	-- LDA @5                      	--Carrega o valor do endereço 5 da RAM no acumulador (Limite das centenas de milhares)
tmp(67) := STA & '1' & x"25";	-- STA @293                    	--Mostra o valor do acumulador HEX 5 (centenas de milhares)
tmp(68) := NOP & '0' & x"00";	-- !LimUni
tmp(69) := LDA & '1' & x"40";	-- LDA @320                    	--Carrega valor das chaves SW0 a SW7 no acumulador
tmp(70) := CEQ & '0' & x"14";	-- CEQ @20                     	--Compara o valor das chaves SW0 a SW7 com 20 (10)
tmp(71) := JEQ & '0' & x"55";	-- JEQ @maxUni                 	--Se o valor das chaves SW0 a SW7 for 10, vai para o label maxUni (Limite maximo das unidades)
tmp(72) := CEQ & '0' & x"15";	-- CEQ @21                     	--Compara o valor das chaves SW0 a SW7 com 21 (11)
tmp(73) := JEQ & '0' & x"55";	-- JEQ @maxUni                 	--Se o valor das chaves SW0 a SW7 for 11, vai para o label maxUni (Limite maximo das unidades)
tmp(74) := CEQ & '0' & x"16";	-- CEQ @22                     	--Compara o valor das chaves SW0 a SW7 com 22 (12)
tmp(75) := JEQ & '0' & x"55";	-- JEQ @maxUni                 	--Se o valor das chaves SW0 a SW7 for 12, vai para o label maxUni (Limite maximo das unidades)
tmp(76) := CEQ & '0' & x"17";	-- CEQ @23                     	--Compara o valor das chaves SW0 a SW7 com 23 (13)
tmp(77) := JEQ & '0' & x"55";	-- JEQ @maxUni                 	--Se o valor das chaves SW0 a SW7 for 13, vai para o label maxUni (Limite maximo das unidades)
tmp(78) := CEQ & '0' & x"18";	-- CEQ @24                     	--Compara o valor das chaves SW0 a SW7 com 24 (14)
tmp(79) := JEQ & '0' & x"55";	-- JEQ @maxUni                 	--Se o valor das chaves SW0 a SW7 for 14, vai para o label maxUni (Limite maximo das unidades)
tmp(80) := CEQ & '0' & x"19";	-- CEQ @25                     	--Compara o valor das chaves SW0 a SW7 com 25 (15)
tmp(81) := JEQ & '0' & x"55";	-- JEQ @maxUni                 	--Se o valor das chaves SW0 a SW7 for 15, vai para o label maxUni (Limite maximo das unidades)
tmp(82) := STA & '1' & x"20";	-- STA @288                    	--Mostra o valor do acumulador HEX 0 (unidades)
tmp(83) := STA & '0' & x"00";	-- STA @0                      	--Salva o valor do acumulador no endereço 0 da RAM (Limite das unidades)
tmp(84) := JMP & '0' & x"59";	-- JMP @UNIOK                  	--Vai para o label UNIOK (Unidades menor que o limite)
tmp(85) := NOP & '0' & x"00";	-- !maxUni
tmp(86) := LDA & '0' & x"13";	-- LDA @19                     	--Carrega o endereco 19 da RAM no acumulador (9)
tmp(87) := STA & '1' & x"20";	-- STA @288                    	--Mostra o valor do acumulador HEX 0 (unidades)
tmp(88) := STA & '0' & x"00";	-- STA @0                      	--Salva 9 no endereço 0 da RAM (Limite das unidades)
tmp(89) := NOP & '0' & x"00";	-- !UNIOK
tmp(90) := LDA & '1' & x"61";	-- LDA @353                    	--Carrega o valor do KEY1 no acumulador
tmp(91) := CEQ & '0' & x"3E";	-- CEQ @62                     	--Compara o valor do KEY1 com 62 (0)
tmp(92) := JEQ & '0' & x"44";	-- JEQ @LimUni                 	--Se o valor do KEY1 for 0 (nao setou o limite das unidades), vai para o label LimUni (Limite das unidades)
tmp(93) := STA & '1' & x"FE";	-- STA @510                    	--Limpa leitura KEY1
tmp(94) := NOP & '0' & x"00";	-- !LimDez
tmp(95) := LDA & '1' & x"40";	-- LDA @320                    	--Carrega valor das chaves SW0 a SW7 no acumulador
tmp(96) := CEQ & '0' & x"14";	-- CEQ @20                     	--Compara o valor das chaves SW0 a SW7 com 20 (10)
tmp(97) := JEQ & '0' & x"6F";	-- JEQ @maxDez                 	--Se o valor das chaves SW0 a SW7 for 10, vai para o label maxDez (Limite maximo das dezenas)
tmp(98) := CEQ & '0' & x"15";	-- CEQ @21                     	--Compara o valor das chaves SW0 a SW7 com 21 (11)
tmp(99) := JEQ & '0' & x"6F";	-- JEQ @maxDez                 	--Se o valor das chaves SW0 a SW7 for 11, vai para o label maxDez (Limite maximo das dezenas)
tmp(100) := CEQ & '0' & x"16";	-- CEQ @22                     	--Compara o valor das chaves SW0 a SW7 com 22 (12)
tmp(101) := JEQ & '0' & x"6F";	-- JEQ @maxDez                 	--Se o valor das chaves SW0 a SW7 for 12, vai para o label maxDez (Limite maximo das dezenas)
tmp(102) := CEQ & '0' & x"17";	-- CEQ @23                     	--Compara o valor das chaves SW0 a SW7 com 23 (13)
tmp(103) := JEQ & '0' & x"6F";	-- JEQ @maxDez                 	--Se o valor das chaves SW0 a SW7 for 13, vai para o label maxDez (Limite maximo das dezenas)
tmp(104) := CEQ & '0' & x"18";	-- CEQ @24                     	--Compara o valor das chaves SW0 a SW7 com 24 (14)
tmp(105) := JEQ & '0' & x"6F";	-- JEQ @maxDez                 	--Se o valor das chaves SW0 a SW7 for 14, vai para o label maxDez (Limite maximo das dezenas)
tmp(106) := CEQ & '0' & x"19";	-- CEQ @25                     	--Compara o valor das chaves SW0 a SW7 com 25 (15)
tmp(107) := JEQ & '0' & x"6F";	-- JEQ @maxDez                 	--Se o valor das chaves SW0 a SW7 for 15, vai para o label maxDez (Limite maximo das dezenas)
tmp(108) := STA & '1' & x"21";	-- STA @289                    	--Mostra o valor do acumulador HEX 1 (dezenas)
tmp(109) := STA & '0' & x"01";	-- STA @1                      	--Salva o valor do acumulador no endereço 1 da RAM (Limite das dezenas)
tmp(110) := JMP & '0' & x"73";	-- JMP @DEZOK                  	--Vai para o label DEZOK (Dezenas menor que o limite)
tmp(111) := NOP & '0' & x"00";	-- !maxDez
tmp(112) := LDA & '0' & x"13";	-- LDA @19                     	--Carrega 19 no acumulador
tmp(113) := STA & '1' & x"21";	-- STA @289                    	--Mostra o valor do acumulador HEX 1 (dezenas)
tmp(114) := STA & '0' & x"01";	-- STA @1                      	--Salva 9 no endereço 1 da RAM (Limite das dezenas)
tmp(115) := NOP & '0' & x"00";	-- !DEZOK
tmp(116) := LDA & '1' & x"61";	-- LDA @353                    	--Carrega o valor do KEY1 no acumulador
tmp(117) := CEQ & '0' & x"3E";	-- CEQ @62                     	--Compara o valor do KEY1 com 62 (0)
tmp(118) := JEQ & '0' & x"5E";	-- JEQ @LimDez                 	--Se o valor do KEY1 for 0 (nao setou o limite das dezenas), vai para o label LimDez (Limite das dezenas)
tmp(119) := STA & '1' & x"FE";	-- STA @510                    	--Limpa leitura KEY1
tmp(120) := NOP & '0' & x"00";	-- !LimCen
tmp(121) := LDA & '1' & x"40";	-- LDA @320                    	--Carrega valor das chaves SW0 a SW7 no acumulador
tmp(122) := CEQ & '0' & x"14";	-- CEQ @20                     	--Compara o valor das chaves SW0 a SW7 com 20 (10)
tmp(123) := JEQ & '0' & x"89";	-- JEQ @maxCen                 	--Se o valor das chaves SW0 a SW7 for 10, vai para o label maxCen (Limite maximo das centenas)
tmp(124) := CEQ & '0' & x"15";	-- CEQ @21                     	--Compara o valor das chaves SW0 a SW7 com 21 (11)
tmp(125) := JEQ & '0' & x"89";	-- JEQ @maxCen                 	--Se o valor das chaves SW0 a SW7 for 11, vai para o label maxCen (Limite maximo das centenas)
tmp(126) := CEQ & '0' & x"16";	-- CEQ @22                     	--Compara o valor das chaves SW0 a SW7 com 22 (12)
tmp(127) := JEQ & '0' & x"89";	-- JEQ @maxCen                 	--Se o valor das chaves SW0 a SW7 for 12, vai para o label maxCen (Limite maximo das centenas)
tmp(128) := CEQ & '0' & x"17";	-- CEQ @23                     	--Compara o valor das chaves SW0 a SW7 com 23 (13)
tmp(129) := JEQ & '0' & x"89";	-- JEQ @maxCen                 	--Se o valor das chaves SW0 a SW7 for 13, vai para o label maxCen (Limite maximo das centenas)
tmp(130) := CEQ & '0' & x"18";	-- CEQ @24                     	--Compara o valor das chaves SW0 a SW7 com 24 (14)
tmp(131) := JEQ & '0' & x"89";	-- JEQ @maxCen                 	--Se o valor das chaves SW0 a SW7 for 14, vai para o label maxCen (Limite maximo das centenas)
tmp(132) := CEQ & '0' & x"19";	-- CEQ @25                     	--Compara o valor das chaves SW0 a SW7 com 25 (15)
tmp(133) := JEQ & '0' & x"89";	-- JEQ @maxCen                 	--Se o valor das chaves SW0 a SW7 for 15, vai para o label maxCen (Limite maximo das centenas)
tmp(134) := STA & '1' & x"22";	-- STA @290                    	--Mostra o valor do acumulador HEX 2 (centenas)
tmp(135) := STA & '0' & x"02";	-- STA @2                      	--Salva o valor do acumulador no endereço 2 da RAM (Limite das centenas)
tmp(136) := JMP & '0' & x"8D";	-- JMP @CENOK                  	--Vai para o label CENOK (Centenas menor que o limite)
tmp(137) := NOP & '0' & x"00";	-- !maxCen
tmp(138) := LDA & '0' & x"13";	-- LDA @19                     	--Carrega 19 no acumulador
tmp(139) := STA & '1' & x"22";	-- STA @290                    	--Mostra o valor do acumulador HEX 2 (centenas)
tmp(140) := STA & '0' & x"02";	-- STA @2                      	--Salva 9 no endereço 2 da RAM (Limite das centenas)
tmp(141) := NOP & '0' & x"00";	-- !CENOK
tmp(142) := LDA & '1' & x"61";	-- LDA @353                    	--Carrega o valor do KEY1 no acumulador
tmp(143) := CEQ & '0' & x"3E";	-- CEQ @62                     	--Compara o valor do KEY1 com 62 (0)
tmp(144) := JEQ & '0' & x"78";	-- JEQ @LimCen                 	--Se o valor do KEY1 for 0 (nao setou o limite das centenas), vai para o label LimCen (Limite das centenas)
tmp(145) := STA & '1' & x"FE";	-- STA @510                    	--Limpa leitura KEY1
tmp(146) := NOP & '0' & x"00";	-- !LimMil
tmp(147) := LDA & '1' & x"40";	-- LDA @320                    	--Carrega valor das chaves SW0 a SW7 no acumulador
tmp(148) := CEQ & '0' & x"14";	-- CEQ @20                     	--Compara o valor das chaves SW0 a SW7 com 20 (10)
tmp(149) := JEQ & '0' & x"A3";	-- JEQ @maxMil                 	--Se o valor das chaves SW0 a SW7 for 10, vai para o label maxMil (Limite maximo dos milhares)
tmp(150) := CEQ & '0' & x"15";	-- CEQ @21                     	--Compara o valor das chaves SW0 a SW7 com 21 (11)
tmp(151) := JEQ & '0' & x"A3";	-- JEQ @maxMil                 	--Se o valor das chaves SW0 a SW7 for 11, vai para o label maxMil (Limite maximo dos milhares)
tmp(152) := CEQ & '0' & x"16";	-- CEQ @22                     	--Compara o valor das chaves SW0 a SW7 com 22 (12)
tmp(153) := JEQ & '0' & x"A3";	-- JEQ @maxMil                 	--Se o valor das chaves SW0 a SW7 for 12, vai para o label maxMil (Limite maximo dos milhares)
tmp(154) := CEQ & '0' & x"17";	-- CEQ @23                     	--Compara o valor das chaves SW0 a SW7 com 23 (13)
tmp(155) := JEQ & '0' & x"A3";	-- JEQ @maxMil                 	--Se o valor das chaves SW0 a SW7 for 13, vai para o label maxMil (Limite maximo dos milhares)
tmp(156) := CEQ & '0' & x"18";	-- CEQ @24                     	--Compara o valor das chaves SW0 a SW7 com 24 (14)
tmp(157) := JEQ & '0' & x"A3";	-- JEQ @maxMil                 	--Se o valor das chaves SW0 a SW7 for 14, vai para o label maxMil (Limite maximo dos milhares)
tmp(158) := CEQ & '0' & x"19";	-- CEQ @25                     	--Compara o valor das chaves SW0 a SW7 com 25 (15)
tmp(159) := JEQ & '0' & x"A3";	-- JEQ @maxMil                 	--Se o valor das chaves SW0 a SW7 for 15, vai para o label maxMil (Limite maximo dos milhares)
tmp(160) := STA & '1' & x"23";	-- STA @291                    	--Mostra o valor do acumulador HEX 3 (milhares)
tmp(161) := STA & '0' & x"03";	-- STA @3                      	--Salva o valor do acumulador no endereço 3 da RAM (Limite dos milhares)
tmp(162) := JMP & '0' & x"A7";	-- JMP @MILOK                  	--Vai para o label MILOK (Milhares menor que o limite)
tmp(163) := NOP & '0' & x"00";	-- !maxMil
tmp(164) := LDA & '0' & x"13";	-- LDA @19                     	--Carrega 19 no acumulador
tmp(165) := STA & '1' & x"23";	-- STA @291                    	--Mostra o valor do acumulador HEX 3 (milhares)
tmp(166) := STA & '0' & x"03";	-- STA @3                      	--Salva 9 no endereço 3 da RAM (Limite dos milhares)
tmp(167) := NOP & '0' & x"00";	-- !MILOK
tmp(168) := LDA & '1' & x"61";	-- LDA @353                    	--Carrega o valor do KEY1 no acumulador
tmp(169) := CEQ & '0' & x"3E";	-- CEQ @62                     	--Compara o valor do KEY1 com 62 (0)
tmp(170) := JEQ & '0' & x"92";	-- JEQ @LimMil                 	--Se o valor do KEY1 for 0 (nao setou o limite dos milhares), vai para o label LimMil (Limite dos milhares)
tmp(171) := STA & '1' & x"FE";	-- STA @510                    	--Limpa leitura KEY1
tmp(172) := NOP & '0' & x"00";	-- !LimDezM
tmp(173) := LDA & '1' & x"40";	-- LDA @320                    	--Carrega valor das chaves SW0 a SW7 no acumulador
tmp(174) := CEQ & '0' & x"14";	-- CEQ @20                     	--Compara o valor das chaves SW0 a SW7 com 20 (10)
tmp(175) := JEQ & '0' & x"6F";	-- JEQ @maxDezM                	--Se o valor das chaves SW0 a SW7 for 10, vai para o label maxDezM (Limite maximo das dezenas de milhares)
tmp(176) := CEQ & '0' & x"15";	-- CEQ @21                     	--Compara o valor das chaves SW0 a SW7 com 21 (11)
tmp(177) := JEQ & '0' & x"6F";	-- JEQ @maxDezM                	--Se o valor das chaves SW0 a SW7 for 11, vai para o label maxDezM (Limite maximo das dezenas de milhares)
tmp(178) := CEQ & '0' & x"16";	-- CEQ @22                     	--Compara o valor das chaves SW0 a SW7 com 22 (12)
tmp(179) := JEQ & '0' & x"6F";	-- JEQ @maxDezM                	--Se o valor das chaves SW0 a SW7 for 12, vai para o label maxDezM (Limite maximo das dezenas de milhares)
tmp(180) := CEQ & '0' & x"17";	-- CEQ @23                     	--Compara o valor das chaves SW0 a SW7 com 23 (13)
tmp(181) := JEQ & '0' & x"6F";	-- JEQ @maxDezM                	--Se o valor das chaves SW0 a SW7 for 13, vai para o label maxDezM (Limite maximo das dezenas de milhares)
tmp(182) := CEQ & '0' & x"18";	-- CEQ @24                     	--Compara o valor das chaves SW0 a SW7 com 24 (14)
tmp(183) := JEQ & '0' & x"6F";	-- JEQ @maxDezM                	--Se o valor das chaves SW0 a SW7 for 14, vai para o label maxDezM (Limite maximo das dezenas de milhares)
tmp(184) := CEQ & '0' & x"19";	-- CEQ @25                     	--Compara o valor das chaves SW0 a SW7 com 25 (15)
tmp(185) := JEQ & '0' & x"6F";	-- JEQ @maxDezM                	--Se o valor das chaves SW0 a SW7 for 15, vai para o label maxDezM (Limite maximo das dezenas de milhares)
tmp(186) := STA & '1' & x"24";	-- STA @292                    	--Mostra o valor do acumulador HEX 4 (dezenas de milhares)
tmp(187) := STA & '0' & x"04";	-- STA @4                      	--Salva o valor do acumulador no endereço 4 da RAM (Limite das dezenas de milhares)
tmp(188) := JMP & '0' & x"C1";	-- JMP @DEZMOK                 	--Vai para o label DEZMOK (Dezenas de milhares menor que o limite)
tmp(189) := NOP & '0' & x"00";	-- !maxDezM
tmp(190) := LDA & '0' & x"13";	-- LDA @19                     	--Carrega 19 no acumulador
tmp(191) := STA & '1' & x"24";	-- STA @292                    	--Mostra o valor do acumulador HEX 4 (dezenas de milhares)
tmp(192) := STA & '0' & x"04";	-- STA @4                      	--Salva 9 no endereço 4 da RAM (Limite das dezenas de milhares)
tmp(193) := NOP & '0' & x"00";	-- !DEZMOK
tmp(194) := LDA & '1' & x"61";	-- LDA @353                    	--Carrega o valor do KEY1 no acumulador
tmp(195) := CEQ & '0' & x"3E";	-- CEQ @62                     	--Compara o valor do KEY1 com 62 (0)
tmp(196) := JEQ & '0' & x"5E";	-- JEQ @LimDezM                	--Se o valor do KEY1 for 0 (nao setou o limite das dezenas de milhares), vai para o label LimDezM (Limite das dezenas de milhares)
tmp(197) := STA & '1' & x"FE";	-- STA @510                    	--Limpa leitura KEY1
tmp(198) := NOP & '0' & x"00";	-- !LimCenM
tmp(199) := LDA & '1' & x"40";	-- LDA @320                    	--Carrega valor das chaves SW0 a SW7 no acumulador
tmp(200) := CEQ & '0' & x"14";	-- CEQ @20                     	--Compara o valor das chaves SW0 a SW7 com 20 (10)
tmp(201) := JEQ & '0' & x"89";	-- JEQ @maxCenM                	--Se o valor das chaves SW0 a SW7 for 10, vai para o label maxCenM (Limite maximo das centenas de milhares)
tmp(202) := CEQ & '0' & x"15";	-- CEQ @21                     	--Compara o valor das chaves SW0 a SW7 com 21 (11)
tmp(203) := JEQ & '0' & x"89";	-- JEQ @maxCenM                	--Se o valor das chaves SW0 a SW7 for 11, vai para o label maxCenM (Limite maximo das centenas de milhares)
tmp(204) := CEQ & '0' & x"16";	-- CEQ @22                     	--Compara o valor das chaves SW0 a SW7 com 22 (12)
tmp(205) := JEQ & '0' & x"89";	-- JEQ @maxCenM                	--Se o valor das chaves SW0 a SW7 for 12, vai para o label maxCenM (Limite maximo das centenas de milhares)
tmp(206) := CEQ & '0' & x"17";	-- CEQ @23                     	--Compara o valor das chaves SW0 a SW7 com 23 (13)
tmp(207) := JEQ & '0' & x"89";	-- JEQ @maxCenM                	--Se o valor das chaves SW0 a SW7 for 13, vai para o label maxCenM (Limite maximo das centenas de milhares)
tmp(208) := CEQ & '0' & x"18";	-- CEQ @24                     	--Compara o valor das chaves SW0 a SW7 com 24 (14)
tmp(209) := JEQ & '0' & x"89";	-- JEQ @maxCenM                	--Se o valor das chaves SW0 a SW7 for 14, vai para o label maxCenM (Limite maximo das centenas de milhares)
tmp(210) := CEQ & '0' & x"19";	-- CEQ @25                     	--Compara o valor das chaves SW0 a SW7 com 25 (15)
tmp(211) := JEQ & '0' & x"89";	-- JEQ @maxCenM                	--Se o valor das chaves SW0 a SW7 for 15, vai para o label maxCenM (Limite maximo das centenas de milhares)
tmp(212) := STA & '1' & x"25";	-- STA @293                    	--Mostra o valor do acumulador HEX 5 (centenas de milhares)
tmp(213) := STA & '0' & x"05";	-- STA @5                      	--Salva o valor do acumulador no endereço 5 da RAM (Limite das centenas de milhares)
tmp(214) := JMP & '0' & x"DB";	-- JMP @CENMOK                 	--Vai para o label CENMOK (Centenas de milhares menor que o limite)
tmp(215) := NOP & '0' & x"00";	-- !maxCenM
tmp(216) := LDA & '0' & x"13";	-- LDA @19                     	--Carrega 19 no acumulador
tmp(217) := STA & '1' & x"25";	-- STA @293                    	--Mostra o valor do acumulador HEX 5 (centenas de milhares)
tmp(218) := STA & '0' & x"05";	-- STA @5                      	--Salva 9 no endereço 5 da RAM (Limite das centenas de milhares)
tmp(219) := NOP & '0' & x"00";	-- !CENMOK
tmp(220) := LDA & '1' & x"61";	-- LDA @353                    	--Carrega o valor do KEY1 no acumulador
tmp(221) := CEQ & '0' & x"3E";	-- CEQ @62                     	--Compara o valor do KEY1 com 62 (0)
tmp(222) := JEQ & '0' & x"78";	-- JEQ @LimCenM                	--Se o valor do KEY1 for 0 (nao setou o limite das centenas de milhares), vai para o label LimCenM (Limite das centenas de milhares)
tmp(223) := STA & '1' & x"FE";	-- STA @510                    	--Limpa leitura KEY1
tmp(224) := LDA & '0' & x"0A";	-- LDA @10                     	--Carrega o valor do endereço 10 da RAM no acumulador (valor atual das unidades)
tmp(225) := STA & '1' & x"20";	-- STA @288                    	--Mostra o valor do acumulador HEX 0 (unidades)
tmp(226) := LDA & '0' & x"0B";	-- LDA @11                     	--Carrega o valor do endereço 11 da RAM no acumulador (valor atual das dezenas)
tmp(227) := STA & '1' & x"21";	-- STA @289                    	--Mostra o valor do acumulador HEX 1 (dezenas)
tmp(228) := LDA & '0' & x"0C";	-- LDA @12                     	--Carrega o valor do endereço 12 da RAM no acumulador (valor atual das centenas)
tmp(229) := STA & '1' & x"22";	-- STA @290                    	--Mostra o valor do acumulador HEX 2 (centenas)
tmp(230) := LDA & '0' & x"0D";	-- LDA @13                     	--Carrega o valor do endereço 13 da RAM no acumulador (valor atual dos milhares)
tmp(231) := STA & '1' & x"23";	-- STA @291                    	--Mostra o valor do acumulador HEX 3 (milhares)
tmp(232) := LDA & '0' & x"0E";	-- LDA @14                     	--Carrega o valor do endereço 14 da RAM no acumulador (valor atual das dezenas de milhares)
tmp(233) := STA & '1' & x"24";	-- STA @292                    	--Mostra o valor do acumulador HEX 4 (dezenas de milhares)
tmp(234) := LDA & '0' & x"0F";	-- LDA @15                     	--Carrega o valor do endereço 15 da RAM no acumulador (valor atual das centenas de milhares)
tmp(235) := STA & '1' & x"25";	-- STA @293                    	--Mostra o valor do acumulador HEX 5 (centenas de milhares)
tmp(236) := JMP & '0' & x"2B";	-- JMP @Start                  	--Volta para o label Start (inicio do programa)
tmp(237) := NOP & '0' & x"00";	-- !Incremento
tmp(238) := STA & '1' & x"FF";	-- STA @511                    	--Limpa leitura KEY0
tmp(239) := LDA & '0' & x"0A";	-- LDA @10                     	--Carrega o valor do endereço 10 da RAM no acumulador (valor atual das unidades)
tmp(240) := SOMA & '0' & x"3F";	-- SOMA @63                    	--Soma o valor do acumulador com 63 (1)
tmp(241) := CEQ & '0' & x"14";	-- CEQ @20                     	--Compara o valor do acumulador com o endereco 20 da RAM (10)
tmp(242) := JEQ & '0' & x"F5";	-- JEQ @IncDez                 	--Se o valor do acumulador for 10, vai para o label IncDez (Incremento das dezenas)
tmp(243) := STA & '0' & x"0A";	-- STA @10                     	--Se o valor do acumulador nao for 10, salva o valor do acumulador no endereço 10 da RAM (valor atual das unidades)
tmp(244) := JMP & '1' & x"22";	-- JMP @Display                	--Vai para o label Display (Mostra o valor atual)
tmp(245) := NOP & '0' & x"00";	-- !IncDez
tmp(246) := LDA & '0' & x"3E";	-- LDA @62                     	--Carrega o valor 62 (0) no acumulador
tmp(247) := STA & '0' & x"0A";	-- STA @10                     	--Zera o valor atual das unidades
tmp(248) := LDA & '0' & x"0B";	-- LDA @11                     	--Carrega o valor do endereço 11 da RAM no acumulador (valor atual das dezenas)
tmp(249) := SOMA & '0' & x"3F";	-- SOMA @63                    	--Soma o valor do acumulador com 63 (1)
tmp(250) := CEQ & '0' & x"14";	-- CEQ @20                     	--Compara o valor do acumulador com o endereco 20 da RAM (10)
tmp(251) := JEQ & '0' & x"FE";	-- JEQ @IncCen                 	--Se o valor do acumulador for 10, vai para o label IncCen (Incremento das centenas)
tmp(252) := STA & '0' & x"0B";	-- STA @11                     	--Se o valor do acumulador nao for 10, salva o valor do acumulador no endereço 11 da RAM (valor atual das dezenas)
tmp(253) := JMP & '1' & x"22";	-- JMP @Display                	--Vai para o label Display (Mostra o valor atual)
tmp(254) := NOP & '0' & x"00";	-- !IncCen
tmp(255) := LDA & '0' & x"3E";	-- LDA @62                     	--Carrega o valor 62 (0) no acumulador
tmp(256) := STA & '0' & x"0B";	-- STA @11                     	--Zera o valor atual das dezenas
tmp(257) := LDA & '0' & x"0C";	-- LDA @12                     	--Carrega o valor do endereço 12 da RAM no acumulador (valor atual das centenas)
tmp(258) := SOMA & '0' & x"3F";	-- SOMA @63                    	--Soma o valor do acumulador com 63 (1)
tmp(259) := CEQ & '0' & x"14";	-- CEQ @20                     	--Compara o valor do acumulador com o endereco 20 da RAM (10)
tmp(260) := JEQ & '1' & x"07";	-- JEQ @IncMil                 	--Se o valor do acumulador for 10, vai para o label IncMil (Incremento dos milhares)
tmp(261) := STA & '0' & x"0C";	-- STA @12                     	--Se o valor do acumulador nao for 10, salva o valor do acumulador no endereço 12 da RAM (valor atual das centenas)
tmp(262) := JMP & '1' & x"22";	-- JMP @Display                	--Vai para o label Display (Mostra o valor atual)
tmp(263) := NOP & '0' & x"00";	-- !IncMil
tmp(264) := LDA & '0' & x"3E";	-- LDA @62                     	--Carrega o valor 62 (0) no acumulador
tmp(265) := STA & '0' & x"0C";	-- STA @12                     	--Zera o valor atual das centenas
tmp(266) := LDA & '0' & x"0D";	-- LDA @13                     	--Carrega o valor do endereço 13 da RAM no acumulador (valor atual dos milhares)
tmp(267) := SOMA & '0' & x"3F";	-- SOMA @63                    	--Soma o valor do acumulador com 63 (1)
tmp(268) := CEQ & '0' & x"14";	-- CEQ @20                     	--Compara o valor do acumulador com o endereco 20 da RAM (10)
tmp(269) := JEQ & '0' & x"F5";	-- JEQ @IncDezM                	--Se o valor do acumulador for 10, vai para o label IncDezM (Incremento das dezenas de milhares)
tmp(270) := STA & '0' & x"0D";	-- STA @13                     	--Se o valor do acumulador nao for 10, salva o valor do acumulador no endereço 13 da RAM (valor atual dos milhares)
tmp(271) := JMP & '1' & x"22";	-- JMP @Display                	--Vai para o label Display (Mostra o valor atual)
tmp(272) := NOP & '0' & x"00";	-- !IncDezM
tmp(273) := LDA & '0' & x"3E";	-- LDA @62                     	--Carrega o valor 62 (0) no acumulador
tmp(274) := STA & '0' & x"0D";	-- STA @13                     	--Zera o valor atual dos milhares
tmp(275) := LDA & '0' & x"0E";	-- LDA @14                     	--Carrega o valor do endereço 14 da RAM no acumulador (valor atual das dezenas de milhares)
tmp(276) := SOMA & '0' & x"3F";	-- SOMA @63                    	--Soma o valor do acumulador com 63 (1)
tmp(277) := CEQ & '0' & x"14";	-- CEQ @20                     	--Compara o valor do acumulador com o endereco 20 da RAM (10)
tmp(278) := JEQ & '0' & x"FE";	-- JEQ @IncCenM                	--Se o valor do acumulador for 10, vai para o label IncCenM (Incremento das centenas de milhares)
tmp(279) := STA & '0' & x"0E";	-- STA @14                     	--Se o valor do acumulador nao for 10, salva o valor do acumulador no endereço 14 da RAM (valor atual das dezenas de milhares)
tmp(280) := JMP & '1' & x"22";	-- JMP @Display                	--Vai para o label Display (Mostra o valor atual)
tmp(281) := NOP & '0' & x"00";	-- !IncCenM
tmp(282) := LDA & '0' & x"3E";	-- LDA @62                     	--Carrega o valor 62 (0) no acumulador
tmp(283) := STA & '0' & x"0E";	-- STA @14                     	--Zera o valor atual das dezenas de milhares
tmp(284) := LDA & '0' & x"0F";	-- LDA @15                     	--Carrega o valor do endereço 15 da RAM no acumulador (valor atual das centenas de milhares)
tmp(285) := SOMA & '0' & x"3F";	-- SOMA @63                    	--Soma o valor do acumulador com 63 (1)
tmp(286) := CEQ & '0' & x"14";	-- CEQ @20                     	--Compara o valor do acumulador com o endereco 20 da RAM (10)
tmp(287) := JEQ & '1' & x"30";	-- JEQ @NoveNove               	--Se o valor do acumulador for 10, vai para o label NoveNove (valor nos displays igual a 999999)
tmp(288) := STA & '0' & x"0F";	-- STA @15                     	--Se o valor do acumulador nao for 10, salva o valor do acumulador no endereço 15 da RAM (valor atual das centenas de milhares)
tmp(289) := JMP & '1' & x"22";	-- JMP @Display                	--Vai para o label Display (Mostra o valor atual)
tmp(290) := NOP & '0' & x"00";	-- !Display
tmp(291) := LDA & '0' & x"0A";	-- LDA @10                     	--Carrega o valor do endereço 10 da RAM no acumulador (valor atual das unidades)
tmp(292) := STA & '1' & x"20";	-- STA @288                    	--Salva o valor do acumulador no HEX 0
tmp(293) := LDA & '0' & x"0B";	-- LDA @11                     	--Carrega o valor do endereço 11 da RAM no acumulador (valor atual das dezenas)
tmp(294) := STA & '1' & x"21";	-- STA @289                    	--Salva o valor do acumulador no HEX 1
tmp(295) := LDA & '0' & x"0C";	-- LDA @12                     	--Carrega o valor do endereço 12 da RAM no acumulador (valor atual das centenas)
tmp(296) := STA & '1' & x"22";	-- STA @290                    	--Salva o valor do acumulador no HEX 2
tmp(297) := LDA & '0' & x"0D";	-- LDA @13                     	--Carrega o valor do endereço 13 da RAM no acumulador (valor atual dos milhares)
tmp(298) := STA & '1' & x"23";	-- STA @291                    	--Salva o valor do acumulador no HEX 3
tmp(299) := LDA & '0' & x"0E";	-- LDA @14                     	--Carrega o valor do endereço 14 da RAM no acumulador (valor atual das dezenas de milhares)
tmp(300) := STA & '1' & x"24";	-- STA @292                    	--Salva o valor do acumulador no HEX 4
tmp(301) := LDA & '0' & x"0F";	-- LDA @15                     	--Carrega o valor do endereço 15 da RAM no acumulador (valor atual das centenas de milhares)
tmp(302) := STA & '1' & x"25";	-- STA @293                    	--Salva o valor do acumulador no HEX 5
tmp(303) := JMP & '1' & x"37";	-- JMP @CompLim                	--Vai para o label CompLim (Compara o valor atual com o valor do limite)
tmp(304) := NOP & '0' & x"00";	-- !NoveNove
tmp(305) := LDA & '0' & x"3F";	-- LDA @63                     	--Carrega o valor 63 (1) no acumulador
tmp(306) := STA & '1' & x"02";	-- STA @258                    	--Ascende o LED 9
tmp(307) := LDA & '1' & x"64";	-- LDA @356                    	--Carrega o valor do Reset no acumulador
tmp(308) := CEQ & '0' & x"3F";	-- CEQ @63                     	--Compara o valor do acumulador com 63 (1)
tmp(309) := JEQ & '0' & x"00";	-- JEQ @Reset                  	--Se o valor do acumulador for 1, vai para o label Reset (Reseta o programa)
tmp(310) := JMP & '1' & x"30";	-- JMP @NoveNove               	--Se o valor do acumulador nao for 1, vai para o label NoveNove
tmp(311) := NOP & '0' & x"00";	-- !CompLim
tmp(312) := LDA & '0' & x"0A";	-- LDA @10                     	--Carrega o valor do endereço 10 da RAM no acumulador (valor atual das unidades)
tmp(313) := CEQ & '0' & x"00";	-- CEQ @0                      	--Compara o valor do acumulador com o endereco 0 da RAM (limite das unidades)
tmp(314) := JEQ & '1' & x"3C";	-- JEQ @CompDez                	--Se for igual, vai para o label CompDez (Compara o valor atual das dezenas com o valor do limite das dezenas)
tmp(315) := JMP & '0' & x"2B";	-- JMP @Start                  	--Se nao for igual, vai para o label Start (Loop principal)
tmp(316) := NOP & '0' & x"00";	-- !CompDez
tmp(317) := LDA & '0' & x"0B";	-- LDA @11                     	--Carrega o valor do endereço 11 da RAM no acumulador (valor atual das dezenas)
tmp(318) := CEQ & '0' & x"01";	-- CEQ @1                      	--Compara o valor do acumulador com o endereco 1 da RAM (limite das dezenas)
tmp(319) := JEQ & '1' & x"41";	-- JEQ @CompCen                	--Se for igual, vai para o label CompCen (Compara o valor atual das centenas com o valor do limite das centenas)
tmp(320) := JMP & '0' & x"2B";	-- JMP @Start                  	--Se nao for igual, vai para o label Start (Loop principal)
tmp(321) := NOP & '0' & x"00";	-- !CompCen
tmp(322) := LDA & '0' & x"0C";	-- LDA @12                     	--Carrega o valor do endereço 12 da RAM no acumulador (valor atual das centenas)
tmp(323) := CEQ & '0' & x"02";	-- CEQ @2                      	--Compara o valor do acumulador com o endereco 2 da RAM (limite das centenas)
tmp(324) := JEQ & '1' & x"46";	-- JEQ @CompMil                	--Se for igual, vai para o label CompMil (Compara o valor atual dos milhares com o valor do limite dos milhares)
tmp(325) := JMP & '0' & x"2B";	-- JMP @Start                  	--Se nao for igual, vai para o label Start (Loop principal)
tmp(326) := NOP & '0' & x"00";	-- !CompMil
tmp(327) := LDA & '0' & x"0D";	-- LDA @13                     	--Carrega o valor do endereço 13 da RAM no acumulador (valor atual dos milhares)
tmp(328) := CEQ & '0' & x"03";	-- CEQ @3                      	--Compara o valor do acumulador com o endereco 3 da RAM (limite dos milhares)
tmp(329) := JEQ & '1' & x"3C";	-- JEQ @CompDezM               	--Se for igual, vai para o label CompDezM (Compara o valor atual das dezenas de milhares com o valor do limite das dezenas de milhares)
tmp(330) := JMP & '0' & x"2B";	-- JMP @Start                  	--Se nao for igual, vai para o label Start (Loop principal)
tmp(331) := NOP & '0' & x"00";	-- !CompDezM
tmp(332) := LDA & '0' & x"0E";	-- LDA @14                     	--Carrega o valor do endereço 14 da RAM no acumulador (valor atual das dezenas de milhares)
tmp(333) := CEQ & '0' & x"04";	-- CEQ @4                      	--Compara o valor do acumulador com o endereco 4 da RAM (limite das dezenas de milhares)
tmp(334) := JEQ & '1' & x"41";	-- JEQ @CompCenM               	--Se for igual, vai para o label CompCenM (Compara o valor atual das centenas de milhares com o valor do limite das centenas de milhares)
tmp(335) := JMP & '0' & x"2B";	-- JMP @Start                  	--Se nao for igual, vai para o label Start (Loop principal)
tmp(336) := NOP & '0' & x"00";	-- !CompCenM
tmp(337) := LDA & '0' & x"0F";	-- LDA @15                     	--Carrega o valor do endereço 15 da RAM no acumulador (valor atual das centenas de milhares)
tmp(338) := CEQ & '0' & x"05";	-- CEQ @5                      	--Compara o valor do acumulador com o endereco 5 da RAM (limite das centenas de milhares)
tmp(339) := JEQ & '1' & x"55";	-- JEQ @Fim                    	--Se for igual, vai para o label Fim (Fim do programa)
tmp(340) := JMP & '0' & x"2B";	-- JMP @Start                  	--Se nao for igual, vai para o label Start (Loop principal)
tmp(341) := NOP & '0' & x"00";	-- !Fim
tmp(342) := LDA & '0' & x"3F";	-- LDA @63                     	--Carrega o valor 63 (1) no acumulador
tmp(343) := STA & '1' & x"02";	-- STA @258                    	--Ascende o LED 9
tmp(344) := STA & '1' & x"01";	-- STA @257                    	--Ascende o LED 8
tmp(345) := LDI & '0' & x"FF";	-- LDI $255                    	--Carrega o valor 255 no acumulador
tmp(346) := STA & '1' & x"00";	-- STA @256                    	--Ascende os LEDs 7 a 0
tmp(347) := LDA & '1' & x"64";	-- LDA @356                    	--Carrega o valor do Reset no acumulador
tmp(348) := CEQ & '0' & x"3F";	-- CEQ @63                     	--Compara o valor do acumulador com 63 (1)
tmp(349) := JEQ & '0' & x"00";	-- JEQ @Reset                  	--Se o valor do acumulador for 1, vai para o label Reset (Reseta o programa)
tmp(350) := JMP & '1' & x"55";	-- JMP @Fim                    	--Se o valor do acumulador nao for 1, vai para o label Fim


        return tmp;
    end initMemory;

    signal memROM : blocoMemoria := initMemory;

begin
    Dado <= memROM (to_integer(unsigned(Endereco)));
end architecture;